package types_pkg;

typedef struct packed {
    logic valid;
    logic sof;
    logic eol;
} flags_t;

endpackage
