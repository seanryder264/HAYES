module frame_reg #(
    // TODO
) (
    // TODO
);
    
    // This block latches the poles and zeroes to set values for a single frame

endmodule