module func_eval  (
    input wire a_re,
    input wire a_im,
    input wire b_re,
    input wire b_im,
);

// Registers that hold the values of 4 poles and 4 zeroes
// Loaded 

    
endmodule