module pixel_generator(
    input           out_stream_aclk,
    input           s_axi_lite_aclk,
    input           axi_resetn,
    input           periph_resetn,

    // Stream output
    output [31:0]   out_stream_tdata,
    output [3:0]    out_stream_tkeep,
    output          out_stream_tlast,
    input           out_stream_tready,
    output          out_stream_tvalid,
    output [0:0]    out_stream_tuser,

    // AXI-Lite S
    input [AXI_LITE_ADDR_WIDTH-1:0]     s_axi_lite_araddr,
    output          s_axi_lite_arready,
    input           s_axi_lite_arvalid,

    input [AXI_LITE_ADDR_WIDTH-1:0]     s_axi_lite_awaddr,
    output          s_axi_lite_awready,
    input           s_axi_lite_awvalid,

    input           s_axi_lite_bready,
    output [1:0]    s_axi_lite_bresp,
    output          s_axi_lite_bvalid,

    output [31:0]   s_axi_lite_rdata,
    input           s_axi_lite_rready,
    output [1:0]    s_axi_lite_rresp,
    output          s_axi_lite_rvalid,

    input  [31:0]   s_axi_lite_wdata,
    output          s_axi_lite_wready,
    input           s_axi_lite_wvalid,

    output [7:0]    r, g, b
);

parameter  REG_FILE_SIZE = 8;
localparam REG_ADDR_WIDTH = $clog2(REG_FILE_SIZE);
localparam REG_FILE_AWIDTH = $clog2(REG_FILE_SIZE);
parameter  AXI_LITE_ADDR_WIDTH = 8;

localparam AWAIT_WADD_AND_DATA = 3'b000;
localparam AWAIT_WDATA = 3'b001;
localparam AWAIT_WADD = 3'b010;
localparam AWAIT_WRITE = 3'b100;
localparam AWAIT_RESP = 3'b101;

localparam AWAIT_RADD = 2'b00;
localparam AWAIT_FETCH = 2'b01;
localparam AWAIT_READ = 2'b10;

localparam AXI_OK = 2'b00;
localparam AXI_ERR = 2'b10;

reg [31:0]                          regfile [REG_FILE_SIZE-1:0];
reg [REG_FILE_AWIDTH-1:0]           writeAddr, readAddr;
reg [31:0]                          readData, writeData;
reg [1:0]                           readState = AWAIT_RADD;
reg [2:0]                           writeState = AWAIT_WADD_AND_DATA;

//Read from the register file
always @(posedge s_axi_lite_aclk) begin
    
    readData <= regfile[readAddr];

    if (!axi_resetn) begin
    readState <= AWAIT_RADD;
    end

    else case (readState)

        AWAIT_RADD: begin
            if (s_axi_lite_arvalid) begin
                readAddr <= s_axi_lite_araddr[2+:REG_FILE_AWIDTH];
                readState <= AWAIT_FETCH;
            end
        end

        AWAIT_FETCH: begin
            readState <= AWAIT_READ;
        end

        AWAIT_READ: begin
            if (s_axi_lite_rready) begin
                readState <= AWAIT_RADD;
            end
        end

        default: begin
            readState <= AWAIT_RADD;
        end

    endcase
end

assign s_axi_lite_arready = (readState == AWAIT_RADD);
assign s_axi_lite_rresp = ({{(REG_ADDR_WIDTH-3){1'b0}}, readAddr} < REG_FILE_SIZE) ? AXI_OK : AXI_ERR;
assign s_axi_lite_rvalid = (readState == AWAIT_READ);
assign s_axi_lite_rdata = readData;

//Write to the register file, use a state machine to track address write, data write and response read events
always @(posedge s_axi_lite_aclk) begin

    if (!axi_resetn) begin
        writeState <= AWAIT_WADD_AND_DATA;
    end

    else case (writeState)

        AWAIT_WADD_AND_DATA: begin  //Idle, awaiting a write address or data
            case ({s_axi_lite_awvalid, s_axi_lite_wvalid})
                2'b10: begin
                    writeAddr <= s_axi_lite_awaddr[2+:REG_FILE_AWIDTH];
                    writeState <= AWAIT_WDATA;
                end
                2'b01: begin
                    writeData <= s_axi_lite_wdata;
                    writeState <= AWAIT_WADD;
                end
                2'b11: begin
                    writeData <= s_axi_lite_wdata;
                    writeAddr <= s_axi_lite_awaddr[2+:REG_FILE_AWIDTH];
                    writeState <= AWAIT_WRITE;
                end
                default: begin
                    writeState <= AWAIT_WADD_AND_DATA;
                end
            endcase        
        end

        AWAIT_WDATA: begin //Received address, waiting for data
            if (s_axi_lite_wvalid) begin
                writeData <= s_axi_lite_wdata;
                writeState <= AWAIT_WRITE;
            end
        end

        AWAIT_WADD: begin //Received data, waiting for address
            if (s_axi_lite_awvalid) begin
                writeAddr <= s_axi_lite_awaddr[2+:REG_FILE_AWIDTH];
                writeState <= AWAIT_WRITE;
            end
        end

        AWAIT_WRITE: begin //Perform the write
            regfile[writeAddr] <= writeData;
            writeState <= AWAIT_RESP;
        end

        AWAIT_RESP: begin //Wait to send response
            if (s_axi_lite_bready) begin
                writeState <= AWAIT_WADD_AND_DATA;
            end
        end

        default: begin
            writeState <= AWAIT_WADD_AND_DATA;
        end
    endcase
end

assign s_axi_lite_awready = (writeState == AWAIT_WADD_AND_DATA || writeState == AWAIT_WADD);
assign s_axi_lite_wready = (writeState == AWAIT_WADD_AND_DATA || writeState == AWAIT_WDATA);
assign s_axi_lite_bvalid = (writeState == AWAIT_RESP);
assign s_axi_lite_bresp = ({{(REG_ADDR_WIDTH-3){1'b0}}, writeAddr} < REG_FILE_SIZE) ? AXI_OK : AXI_ERR;

    wire signed [15:0] x_re;
    wire signed [15:0] y_im;
    wire first, lastx, ready, valid_int;

    // Individual zero/pole registers
    wire [31:0] latched_zeroes_0, latched_zeroes_1, latched_zeroes_2, latched_zeroes_3;
    wire [31:0] latched_poles_0, latched_poles_1, latched_poles_2, latched_poles_3;

    frame_reg frame_reg_inst (
        .clk(out_stream_aclk),
        .reset(!periph_resetn),
        .frame_done(out_stream_tlast),
        .zero_in_0(regfile[0]), .zero_in_1(regfile[1]), 
        .zero_in_2(regfile[2]), .zero_in_3(regfile[3]),
        .pole_in_0(regfile[4]), .pole_in_1(regfile[5]),
        .pole_in_2(regfile[6]), .pole_in_3(regfile[7]),
        .zero_0(latched_zeroes_0), .zero_1(latched_zeroes_1),
        .zero_2(latched_zeroes_2), .zero_3(latched_zeroes_3),
        .pole_0(latched_poles_0), .pole_1(latched_poles_1),
        .pole_2(latched_poles_2), .pole_3(latched_poles_3)
    );

    coord_gen coord_gen_inst(
        .clk(out_stream_aclk),
        .resetn(periph_resetn),
        .ready(ready),
        .x(x_re),
        .y(y_im),
        .first(first),
        .lastx(lastx),
        .valid(valid_int)
    );

    // Complex sub outputs
    wire signed [15:0] zero_diff_re_0, zero_diff_re_1, zero_diff_re_2, zero_diff_re_3;
    wire signed [15:0] zero_diff_im_0, zero_diff_im_1, zero_diff_im_2, zero_diff_im_3;
    wire signed [15:0] pole_diff_re_0, pole_diff_re_1, pole_diff_re_2, pole_diff_re_3;
    wire signed [15:0] pole_diff_im_0, pole_diff_im_1, pole_diff_im_2, pole_diff_im_3;

    complex_sub complex_sub_inst (
        .x(x_re),
        .y(y_im),
        .zero_0(latched_zeroes_0), .zero_1(latched_zeroes_1),
        .zero_2(latched_zeroes_2), .zero_3(latched_zeroes_3),
        .pole_0(latched_poles_0), .pole_1(latched_poles_1),
        .pole_2(latched_poles_2), .pole_3(latched_poles_3),
        .zero_diff_re_0(zero_diff_re_0), .zero_diff_re_1(zero_diff_re_1),
        .zero_diff_re_2(zero_diff_re_2), .zero_diff_re_3(zero_diff_re_3),
        .zero_diff_im_0(zero_diff_im_0), .zero_diff_im_1(zero_diff_im_1),
        .zero_diff_im_2(zero_diff_im_2), .zero_diff_im_3(zero_diff_im_3),
        .pole_diff_re_0(pole_diff_re_0), .pole_diff_re_1(pole_diff_re_1),
        .pole_diff_re_2(pole_diff_re_2), .pole_diff_re_3(pole_diff_re_3),
        .pole_diff_im_0(pole_diff_im_0), .pole_diff_im_1(pole_diff_im_1),
        .pole_diff_im_2(pole_diff_im_2), .pole_diff_im_3(pole_diff_im_3)
    );

    // Pack differences for phase_eval
    wire [63:0] zero_diff_re_packed = {zero_diff_re_3, zero_diff_re_2, zero_diff_re_1, zero_diff_re_0};
    wire [63:0] zero_diff_im_packed = {zero_diff_im_3, zero_diff_im_2, zero_diff_im_1, zero_diff_im_0};
    wire [63:0] pole_diff_re_packed = {pole_diff_re_3, pole_diff_re_2, pole_diff_re_1, pole_diff_re_0};
    wire [63:0] pole_diff_im_packed = {pole_diff_im_3, pole_diff_im_2, pole_diff_im_1, pole_diff_im_0};

    wire [15:0] phase;

    phase_eval phase_eval_inst (
        .zero_diff_re(zero_diff_re_packed),
        .zero_diff_im(zero_diff_im_packed),
        .pole_diff_re(pole_diff_re_packed),
        .pole_diff_im(pole_diff_im_packed),
        .phase_out(phase)
    );

    colour_map colour_map_inst (
        .phase(phase),
        .r(r),
        .g(g),
        .b(b)
    );

    packer pixel_packer(
        .aclk(out_stream_aclk),
        .aresetn(periph_resetn),
        .r(r),
        .g(g),
        .b(b),
        .eol(lastx),
        .in_stream_ready(ready),
        .valid(valid_int),
        .sof(first),
        .out_stream_tdata(out_stream_tdata),
        .out_stream_tkeep(out_stream_tkeep),
        .out_stream_tlast(out_stream_tlast),
        .out_stream_tready(out_stream_tready),
        .out_stream_tvalid(out_stream_tvalid),
        .out_stream_tuser(out_stream_tuser)
    );

endmodule
