module mag_eval (

);

// Also be a log look up for the log magnitude of the function.This way we can also sum the magnitudes of the logs


endmodule
